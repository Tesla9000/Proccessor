// Name: Dev gupta,Pinkesh Mahawar
// Roll No 210318, 210719



module alu_control(input [5:0] opcode, output[5:0] alucontrol);

assign alucontrol=opcode;
endmodule
// Name: Dev gupta,Pinkesh Mahawar
// Roll No 210318, 210719

module shift_left_2(input [31:0] imme,output[6:0] jump);

assign jump= imme<<2;
endmodule
